library verilog;
use verilog.vl_types.all;
entity eittothreeencoder_vlg_vec_tst is
end eittothreeencoder_vlg_vec_tst;
