library verilog;
use verilog.vl_types.all;
entity cnt_60_vlg_vec_tst is
end cnt_60_vlg_vec_tst;
