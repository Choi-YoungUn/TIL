library verilog;
use verilog.vl_types.all;
entity fourbit_addsub_vlg_vec_tst is
end fourbit_addsub_vlg_vec_tst;
