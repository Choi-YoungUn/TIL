library verilog;
use verilog.vl_types.all;
entity ring_counter_vlg_vec_tst is
end ring_counter_vlg_vec_tst;
