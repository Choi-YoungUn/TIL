library verilog;
use verilog.vl_types.all;
entity demux1x8_pack_proce_vlg_vec_tst is
end demux1x8_pack_proce_vlg_vec_tst;
