library verilog;
use verilog.vl_types.all;
entity onebitfullcomparator_vlg_vec_tst is
end onebitfullcomparator_vlg_vec_tst;
