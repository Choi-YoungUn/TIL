library verilog;
use verilog.vl_types.all;
entity onebitfullcomparator_vlg_check_tst is
    port(
        Xo              : in     vl_logic;
        Yo              : in     vl_logic;
        Zo              : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end onebitfullcomparator_vlg_check_tst;
