library verilog;
use verilog.vl_types.all;
entity eitbit_par_register_vlg_vec_tst is
end eitbit_par_register_vlg_vec_tst;
