library verilog;
use verilog.vl_types.all;
entity mux2x1_vlg_check_tst is
    port(
        y               : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end mux2x1_vlg_check_tst;
