library verilog;
use verilog.vl_types.all;
entity myrommemory_vlg_vec_tst is
end myrommemory_vlg_vec_tst;
