library ieee;
use ieee.std_logic_1164.all;

entity D_FF_q is
port (D : in std_logic;
	   clk : in std_logic;
	   clear : in std_logic;
	   Q : out std_logic);
		end D_FF_q;
		
		architecture behav of D_FF_q is
		
		signal temp : std_logic;
		
		begin 
		process(D, clear, clk)
		begin
		if(clear = '1') then
		temp <= '0';
		elsif(clear'event and clear = '0')then
		temp <= '1';
		elsif(clk'event and clk = '1') then
		temp <= D;
		end if;
		end process;
		Q <= temp;
		
		end behav;