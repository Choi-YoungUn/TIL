library verilog;
use verilog.vl_types.all;
entity onebitfullcomparator_vlg_sample_tst is
    port(
        A               : in     vl_logic;
        B               : in     vl_logic;
        Xi              : in     vl_logic;
        Yi              : in     vl_logic;
        Zi              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end onebitfullcomparator_vlg_sample_tst;
