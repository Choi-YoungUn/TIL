library verilog;
use verilog.vl_types.all;
entity sodavending_mechine_vlg_vec_tst is
end sodavending_mechine_vlg_vec_tst;
