library verilog;
use verilog.vl_types.all;
entity DETclock_vlg_vec_tst is
end DETclock_vlg_vec_tst;
